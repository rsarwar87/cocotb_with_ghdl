---------------------------------------------------------------------
--              Standard VITAL_Primitives Package
--    NOTE:     Xilinx Inc is unable to redistribute source code of 
--              Standard VITAL_Primitives Package to our customers 
--              due to IEEE's copyright. 
-- 
--              VHDL source code of Standard VITAL_Primitives Package 
--              can be licensed from IEEE by directly contacting them. 
--              For more information visit ieee's website at 
--              http://stdsbbs.ieee.org 
---------------------------------------------------------------------------
